* source *
VDD vdd 0 1

* input
VA a 0 dc 1
VB b 0 dc 1
VC c 0 dc 1
VD d 0 dc 1


* MOSFET model
.model PMOS PMOS (LEVEL = 1 VTO = -0.5 KP = 50u)
.model NMOS NMOS (LEVEL = 1 VTO = 0.5 KP = 100u)

* A NAND B
Mpa m_mid a vdd vdd PMOS
Mpb m_mid b vdd vdd PMOS

Mna YB a n_mid 0 NMOS
Mnb n_mid b 0 0 NMOS

* C NAND D
Mpc YB c m_mid vdd PMOS
Mpd YB d vdd m_mid PMOS

Mnc YB c n_mid 0 NMOS
Mnd n_mid d 0 0 NMOS

.control

op
print v(YB)

.endc

.end


