* source
VDD vdd 0 1

* input
VA a 0 0
VB b 0 0
VC c 0 0
VD d 0 0

.dc VA 0 1 1 VB 0 1 1 VC 0 1 1 VD 0 1 1
.print dc v(a) v(b) v(c) v(d) v(YB)

* MOSFET model
.model PMOS PMOS (LEVEL = 1 VTO = -0.5 KP = 50u)
.model NMOS NMOS (LEVEL = 1 VTO = 0.5 KP = 100u)

* A NAND B
Mpa m_mid a vdd vdd PMOS
Mpb m_mid b vdd vdd PMOS

Mna YB a n_mid 0 NMOS
Mnb n_mid b 0 0 NMOS

* C NAND D
Mpc YB c m_mid vdd PMOS
Mpd YB d vdd m_mid PMOS

Mnc YB c n_mid 0 NMOS
Mnd n_mid d 0 0 NMOS

.op
.end


